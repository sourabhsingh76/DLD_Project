module BufferBox(G_i_j, P_i_j, G_i_j, P_i_j);
input G_i_j, P_i_j;
output G_i_j, P_i_j;
endmodule